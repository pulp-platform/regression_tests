
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [8:0]  A,
    output logic [63:0] Q
  );

  const logic [63:0] mem[0:1023] = {
    64'h0840006F0880006F,
    64'h07C0006F0800006F,
    64'h0740006F0780006F,
    64'h06C0006F0700006F,
    64'h0640006F0680006F,
    64'h05C0006F0600006F,
    64'h0540006F0580006F,
    64'h04C0006F0500006F,
    64'h0440006F0480006F,
    64'h03C0006F0400006F,
    64'h0340006F0380006F,
    64'h02C0006F0300006F,
    64'h0240006F0280006F,
    64'h01C0006F0200006F,
    64'h0140006F0180006F,
    64'h00C0006F0100006F,
    64'h0000006F4320006F,
    64'h1A10A7B730200073,
    64'h80E7A22304000737,
    64'h0056961380C7A683,
    64'h8247A68300065963,
    64'h80E7A42380E7AA23,
    64'hB7CD105000738082,
    64'h91C7A78397AA6789,
    64'h2023953E6785E7AD,
    64'h07B7200707370005,
    64'h00370793C15C1000,
    64'h07C20085D793C51C,
    64'hE7B3200F083783C1,
    64'hC55C0FF5F5930107,
    64'h0737FFF687938DD9,
    64'hC95C8FD9C90C7047,
    64'hCD1C0785900007B7,
    64'h10C7A0231A1027B7,
    64'hA423475110D7A223,
    64'h46F112A7A02310E7,
    64'h12E7A42312D7A223,
    64'h27831A103737B795,
    64'h8A07280345118A47,
    64'h0034253788A72023,
    64'h079E97AA04950513,
    64'h0207A6230207A423,
    64'h0207AA230207A823,
    64'h0207AE230207AC23,
    64'h242302A801634505,
    64'hCFCCC3D4C39088A7,
    64'hC7984751CF984715,
    64'h8B0553D80007A423,
    64'h880724238082FF75,
    64'h6485C2261141B7CD,
    64'h46C1C42240848613,
    64'hC6064581962A842A,
    64'h40C4A6833F1994A2,
    64'hE69900D7C86347BD,
    64'h01414492442240B2,
    64'h0613660546C18082,
    64'h4422852296224186,
    64'h45C10692449240B2,
    64'h1A10A7B7B5DD0141,
    64'h669180E7A2236711,
    64'hC8631A10A7374781,
    64'h67111A10A7B700A7,
    64'h0073808280E7A423,
    64'h078580D72A231050,
    64'h0A37C4521101B7DD,
    64'h000A0713CA261C00,
    64'hC64EC84ACC226489,
    64'h678594BACE06C256,
    64'hAE2397BA92F4A023,
    64'hA22392B4A22390A4,
    64'hA7831A102AB74007,
    64'hE793892A547D000A,
    64'h67B700FAA0230027,
    64'hC7C0C780C3C01A10,
    64'hCFC0CF80CBC0CB80,
    64'h89AE455143D8D380,
    64'h43D8C3D8F7F77713,
    64'hA78337A5C3D89B75,
    64'h10000793C38D91C4,
    64'h1A1037B700FAA023,
    64'h8887A6238807A423,
    64'h473D8AE7A0234705,
    64'h000A051388E7A223,
    64'h87931C0017B73DCD,
    64'h27B740C7A8830007,
    64'hA783000787931C00,
    64'h65891C0017379207,
    64'h40F006B3FFF78313,
    64'h0537460142070713,
    64'h1563928585931C00,
    64'h660597AA67890316,
    64'h5196061392C7A023,
    64'hAE231A0005B7962A,
    64'h06139337A2239127,
    64'h22E13D8585934006,
    64'h00F56A63FFC72783,
    64'h6963983E00072803,
    64'hB7C1074106050105,
    64'hFF07FBE300B50833,
    64'h8D75951A953E4308,
    64'h5BE81A1047B7B7ED,
    64'h812111410C47A783,
    64'h8163893D4705C606,
    64'h87634709CF8102E7,
    64'h1A10A7B7ED0102E7,
    64'h105000738007A023,
    64'h357545014585BFF5,
    64'hA7B728198105C119,
    64'h00738007A0231A10,
    64'h45054581BFF51050,
    64'hC422C6061141B7DD,
    64'h00F50D634785C226,
    64'hA001CD0D00A7C463,
    64'h479D02F507634795,
    64'h47B7BFCD02F50163,
    64'h1A1044B7DBE81A10,
    64'h74133D05450558E0,
    64'h978240DCD87D1004,
    64'h35B145014585A001,
    64'h3795BFED45054581,
    64'h00C7936387AA962A,
    64'hFFF5C70305858082,
    64'hB7FDFEE78FA30785,
    64'hDA266985D64E7139,
    64'h8493892ACE5ED84A,
    64'hC66ECA666B894189,
    64'hD256D452DC22DE06,
    64'h94CAC86ACC62D05A,
    64'h9BCA99CA4D813369,
    64'h40C9A78301000CB7,
    64'h005007B704FDE363,
    64'hA22307991A1026B7,
    64'h1A1067B7577D0AF6,
    64'hCB98C7D8C798C3D8,
    64'hD398CFD8CF98CBD8,
    64'hC7934149A703429C,
    64'h0006A023C29C1007,
    64'hA783C3D81A1047B7,
    64'hAA03A00197824109,
    64'hAA830004AB030044,
    64'h0D33E40007B70084,
    64'h656344D84C0100FA,
    64'hBF5904C10D8500EC,
    64'h008AF563920BA403,
    64'h86A29871003A8413,
    64'h85DA8652019D7C63,
    64'h9B229A22311D854A,
    64'hB7F90C05408A8AB3,
    64'h3909854A85DA864A,
    64'h3F09855285CA8622,
    64'h011302002117B7D5,
    64'h81320080006F8761,
    64'h3DB1C60611418582,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000};

  logic [10:0] A_Q;

  always_ff @(posedge CLK or negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule