
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [8:0]  A,
    output logic [63:0] Q
  );

  const logic [63:0] mem[0:1023] = {
    64'h0840006F0880006F,
    64'h07C0006F0800006F,
    64'h0740006F0780006F,
    64'h06C0006F0700006F,
    64'h0640006F0680006F,
    64'h05C0006F0600006F,
    64'h0540006F0580006F,
    64'h04C0006F0500006F,
    64'h0440006F0480006F,
    64'h03C0006F0400006F,
    64'h0340006F0380006F,
    64'h02C0006F0300006F,
    64'h0240006F0280006F,
    64'h01C0006F0200006F,
    64'h0140006F0180006F,
    64'h00C0006F0100006F,
    64'h0000006F4EC0006F,
    64'h1A10A7B730200073,
    64'h80E7A22304000737,
    64'h9593421480C78613,
    64'h86930005DC630056,
    64'h8147869342948247,
    64'hC39880878793C298,
    64'hBFF9105000738082,
    64'h91C7A78397AA6789,
    64'h2023953E6785EBAD,
    64'h07B7200707370005,
    64'h00370793C15C1000,
    64'h97B3200F0837C51C,
    64'hB5B30107E7B3DE85,
    64'h87938DD9C55CEE85,
    64'hC90C70470737FFF6,
    64'h900007B7C95C8FD9,
    64'h1A1027B7CD1C0785,
    64'h8713C31010078713,
    64'h10878693C3141047,
    64'h12078693C2984751,
    64'h124786934671C288,
    64'hC39812878793C290,
    64'h05131A103737BF91,
    64'h439C8A4707938A07,
    64'h0513000528034891,
    64'h2023888707138807,
    64'h0513003425370115,
    64'h8513079E97AA0495,
    64'h8513000520230287,
    64'h85130005202302C7,
    64'h8513000520230307,
    64'h8513000520230347,
    64'h8513000520230387,
    64'h2C630005202303C7,
    64'h873EC30845050218,
    64'h8713C31400C7222B,
    64'h87134695C30C01C7,
    64'h00878713C3140187,
    64'h00072023C31446D1,
    64'h3733439802478793,
    64'h20238082FF6DFC17,
    64'hC2261141B7F10007,
    64'hC422408486136485,
    64'h4581962A842A46C1,
    64'hA6833DD194A2C606,
    64'h00D7C86347BD40C4,
    64'h4492442240B2E699,
    64'h660546C180820141,
    64'h8522962241860613,
    64'h0692449240B24422,
    64'hA7B7B555014145C1,
    64'h6691804787131A10,
    64'h470181478793C314,
    64'h1A10A7B700A74863,
    64'h808280E7A4236711,
    64'h0705C39410500073,
    64'h0437CC221101B7E5,
    64'h00040713C4521C00,
    64'hC64EC84ACA266A09,
    64'h67859A3ACE06C256,
    64'h2E2397BA92FA2023,
    64'hA22392BA222390AA,
    64'hA7831A102AB74007,
    64'hC7B3892A54FD000A,
    64'h67B700FAA023C017,
    64'hC304004787131A10,
    64'h8693C28400878693,
    64'h01078693C28400C7,
    64'hC28401478693C284,
    64'h8693C28401878693,
    64'h02078793C28401C7,
    64'h89AE4551431CC384,
    64'h431CC31CC077B7B3,
    64'h37A1C31CC017B7B3,
    64'h0793C79591CA2783,
    64'h37B700FAA0231000,
    64'h2023888787131A10,
    64'hC30488C787130007,
    64'hC3148A0787134685,
    64'hC398473D88478793,
    64'h17B735E100040513,
    64'hA303000787931C00,
    64'h87931C0027B740C7,
    64'h66859207A7830007,
    64'h0633FFF78E136809,
    64'h079341C68E9340F0,
    64'h1C00053745810004,
    64'h9288081342068693,
    64'h97AA678902659563,
    64'h061392C7A0236605,
    64'h1A0005B7962A5196,
    64'h9337A2239127AE23,
    64'h4545859340060613,
    64'h6A6321D7F7032421,
    64'h98BA20D7F88300E5,
    64'h07C1058501156963,
    64'h7BE3010508B3B7C1,
    64'h953A20D7F503FF17,
    64'h47B7B7E58D719572,
    64'h4308074787131A10,
    64'h35338121C6061141,
    64'hA8630C47A783F645,
    64'hE38D0227A0630017,
    64'hC119355945014585,
    64'h1A10A7B7201D8105,
    64'h105000738007A023,
    64'hB7DD45054581BFF5,
    64'hA0231A10A7B7F565,
    64'hBFF5105000738007,
    64'hC226C422C6061141,
    64'hC463478500152C63,
    64'h2963A001CD1500A7,
    64'hBFDD027524630255,
    64'h074787931A1047B7,
    64'h45054004843EC388,
    64'hD8FD1004F4933BFD,
    64'h978243DC1A1047B7,
    64'h3D1145014585A001,
    64'h3785BFED45054581,
    64'h00C59363962E87AA,
    64'h80AB0015C70B8082,
    64'hC2A6715DBFCD00E7,
    64'hDE4E6A0984AADC52,
    64'hD65EC0CA69859A26,
    64'hDA56C4A2C686D462,
    64'hCE6ED06AD266D85A,
    64'h8BB34C013BA98926,
    64'h40CBA783C6520134,
    64'h1A1026B706FC6463,
    64'h0A468713005007B7,
    64'h1A1067B7C31C0799,
    64'hC21800478613577D,
    64'h8613C21800878613,
    64'h01078613C21800C7,
    64'hC21801478613C218,
    64'h8613C21801878613,
    64'h02078793C21801C7,
    64'h414BA703429CC398,
    64'hA023C29C1007C793,
    64'hC3D81A1047B70006,
    64'hA0019782410BA783,
    64'h7A03418787936785,
    64'h41C78793678520F9,
    64'h8793678520F97D83,
    64'h0B3720F97D034207,
    64'h9B6E42498A93E400,
    64'h000AA6839ACA4C81,
    64'h09410C0500DCE563,
    64'h9207A40347B2BFB1,
    64'h003D0413008D7663,
    64'h010007B7C2043433,
    64'h866E00FB7C6386A2,
    64'h9DA23E95852685D2,
    64'h0C85408D0D339A22,
    64'h852685D28626B7D1,
    64'h856E85A686223685,
    64'h02001117B7D53DE1,
    64'h0080006F7BC10113,
    64'hC606114185828132,
    64'h0000000000003D39,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000,
    64'h0000000000000000};

  logic [10:0] A_Q;

  always_ff @(posedge CLK or negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule